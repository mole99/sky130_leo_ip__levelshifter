* NGSPICE file created from sky130_leo_ip__levelshifter_down.ext - technology: sky130A

.subckt sky130_leo_ip__levelshifter_down VDDOUT OUT IN VGND
X0 OUT.t1 a_259_346# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 VDDOUT.t1 IN.t0 a_259_346# VDDOUT.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X2 VDDOUT.t3 a_259_346# OUT.t0 VDDOUT.t2 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X3 a_259_346# IN.t1 VGND.t3 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
R0 VGND.n63 VGND.n52 68735.8
R1 VGND.n52 VGND.n18 25131.8
R2 VGND.n52 VGND.n51 6755.23
R3 VGND.n51 VGND.n50 1593.88
R4 VGND.n48 VGND.n22 1199.38
R5 VGND.n43 VGND.n20 1199.38
R6 VGND.n32 VGND.n25 1199.38
R7 VGND.n28 VGND.n27 1199.38
R8 VGND.n51 VGND.n14 1150.51
R9 VGND.n63 VGND.n53 704.234
R10 VGND.n82 VGND.n81 704.234
R11 VGND.n57 VGND.n13 652.583
R12 VGND.n75 VGND.n7 652.583
R13 VGND.n83 VGND.n5 652.583
R14 VGND.n64 VGND.n15 652.583
R15 VGND.n26 VGND.n18 645.409
R16 VGND.n50 VGND.n19 645.409
R17 VGND.n58 VGND.n57 585
R18 VGND.n59 VGND.n55 585
R19 VGND.n61 VGND.n60 585
R20 VGND.n17 VGND.n16 585
R21 VGND.n65 VGND.n64 585
R22 VGND.n64 VGND.n63 585
R23 VGND.n66 VGND.n15 585
R24 VGND.n53 VGND.n15 585
R25 VGND.n69 VGND.n68 585
R26 VGND.n70 VGND.n69 585
R27 VGND.n4 VGND.n2 585
R28 VGND.n6 VGND.n4 585
R29 VGND.n84 VGND.n83 585
R30 VGND.n83 VGND.n82 585
R31 VGND.n74 VGND.n7 585
R32 VGND.n82 VGND.n7 585
R33 VGND.n73 VGND.n72 585
R34 VGND.n72 VGND.n6 585
R35 VGND.n71 VGND.n12 585
R36 VGND.n71 VGND.n70 585
R37 VGND.n56 VGND.n13 585
R38 VGND.n53 VGND.n13 585
R39 VGND.n76 VGND.n75 585
R40 VGND.n77 VGND.n10 585
R41 VGND.n79 VGND.n78 585
R42 VGND.n11 VGND.n9 585
R43 VGND.n5 VGND.n3 585
R44 VGND.n81 VGND.n5 585
R45 VGND.n38 VGND.n27 585
R46 VGND.n27 VGND.n26 585
R47 VGND.n40 VGND.n39 585
R48 VGND.n41 VGND.n40 585
R49 VGND.n23 VGND.n22 585
R50 VGND.n22 VGND.n19 585
R51 VGND.n48 VGND.n47 585
R52 VGND.n46 VGND.n21 585
R53 VGND.n45 VGND.n20 585
R54 VGND.n50 VGND.n20 585
R55 VGND.n44 VGND.n43 585
R56 VGND.n43 VGND.n19 585
R57 VGND.n42 VGND.n24 585
R58 VGND.n42 VGND.n41 585
R59 VGND.n33 VGND.n25 585
R60 VGND.n26 VGND.n25 585
R61 VGND.n34 VGND.n32 585
R62 VGND.n30 VGND.n29 585
R63 VGND.n37 VGND.n28 585
R64 VGND.n28 VGND.n18 585
R65 VGND.n82 VGND.n6 419.048
R66 VGND.n21 VGND.n20 417.176
R67 VGND.n42 VGND.n25 417.176
R68 VGND.n43 VGND.n42 417.176
R69 VGND.n30 VGND.n28 417.176
R70 VGND.n40 VGND.n27 417.176
R71 VGND.n40 VGND.n22 417.176
R72 VGND.n41 VGND.n19 404.082
R73 VGND.n70 VGND.n14 285.185
R74 VGND.n63 VGND.n54 244.588
R75 VGND.n63 VGND.n62 244.588
R76 VGND.n81 VGND.n8 244.588
R77 VGND.n81 VGND.n80 244.588
R78 VGND.n0 VGND.t1 237.649
R79 VGND.n71 VGND.n13 229.201
R80 VGND.n72 VGND.n71 229.201
R81 VGND.n72 VGND.n7 229.201
R82 VGND.n9 VGND.n5 229.201
R83 VGND.n79 VGND.n10 229.201
R84 VGND.n69 VGND.n15 229.201
R85 VGND.n69 VGND.n4 229.201
R86 VGND.n83 VGND.n4 229.201
R87 VGND.n64 VGND.n17 229.201
R88 VGND.n61 VGND.n55 229.201
R89 VGND.n50 VGND.n49 215.619
R90 VGND.n31 VGND.n18 215.619
R91 VGND.n26 VGND.t0 213.266
R92 VGND.n70 VGND.t2 209.524
R93 VGND.t2 VGND.n6 209.524
R94 VGND.n41 VGND.t0 190.816
R95 VGND.n49 VGND.n48 153.763
R96 VGND.n32 VGND.n31 153.763
R97 VGND.n49 VGND.n21 153.763
R98 VGND.n31 VGND.n30 153.763
R99 VGND.n53 VGND.n14 133.863
R100 VGND.n86 VGND.t3 131.995
R101 VGND.n80 VGND.n79 95.8286
R102 VGND.n75 VGND.n8 95.8286
R103 VGND.n62 VGND.n61 95.8286
R104 VGND.n57 VGND.n54 95.8286
R105 VGND.n55 VGND.n54 95.8286
R106 VGND.n62 VGND.n17 95.8286
R107 VGND.n10 VGND.n8 95.8286
R108 VGND.n80 VGND.n9 95.8286
R109 VGND.n38 VGND.n37 77.9299
R110 VGND.n47 VGND.n23 77.9299
R111 VGND.n45 VGND.n44 77.9299
R112 VGND.n34 VGND.n33 77.9299
R113 VGND.n58 VGND.n56 43.7338
R114 VGND.n76 VGND.n74 43.7338
R115 VGND.n84 VGND.n3 43.7338
R116 VGND.n66 VGND.n65 43.7338
R117 VGND.n39 VGND.n38 27.1064
R118 VGND.n39 VGND.n23 27.1064
R119 VGND.n47 VGND.n46 27.1064
R120 VGND.n46 VGND.n45 27.1064
R121 VGND.n33 VGND.n24 27.1064
R122 VGND.n44 VGND.n24 27.1064
R123 VGND.n34 VGND.n29 27.1064
R124 VGND.n56 VGND.n12 15.3605
R125 VGND.n73 VGND.n12 15.3605
R126 VGND.n74 VGND.n73 15.3605
R127 VGND.n11 VGND.n3 15.3605
R128 VGND.n78 VGND.n11 15.3605
R129 VGND.n78 VGND.n77 15.3605
R130 VGND.n77 VGND.n76 15.3605
R131 VGND.n68 VGND.n2 15.3605
R132 VGND.n84 VGND.n2 15.3605
R133 VGND.n65 VGND.n16 15.3605
R134 VGND.n60 VGND.n16 15.3605
R135 VGND.n60 VGND.n59 15.3605
R136 VGND.n59 VGND.n58 15.3605
R137 VGND.n2 VGND.n1 9.3005
R138 VGND.n85 VGND.n84 9.3005
R139 VGND.n35 VGND.n34 9.3005
R140 VGND.n37 VGND.n36 5.58699
R141 VGND.n36 VGND.n29 5.49833
R142 VGND.n67 VGND.n66 4.25641
R143 VGND.n68 VGND.n67 4.18886
R144 VGND.n67 VGND.n1 2.72752
R145 VGND.n36 VGND.n35 2.06755
R146 VGND.n87 VGND.n86 0.560917
R147 VGND.n35 VGND.n0 0.430708
R148 VGND VGND.n87 0.3385
R149 VGND.n85 VGND.n1 0.1505
R150 VGND.n86 VGND.n85 0.10675
R151 VGND.n87 VGND.n0 0.053
R152 OUT.n0 OUT.t0 356.536
R153 OUT.n0 OUT.t1 237.611
R154 OUT OUT.n0 5.33508
R155 IN.n0 IN.t1 245.971
R156 IN.n0 IN.t0 217.417
R157 IN IN.n0 4.71567
R158 VDDOUT.n27 VDDOUT.n15 681.178
R159 VDDOUT.n21 VDDOUT.n13 681.178
R160 VDDOUT.n38 VDDOUT.n37 681.178
R161 VDDOUT.n35 VDDOUT.n7 681.178
R162 VDDOUT.n82 VDDOUT.t1 663.312
R163 VDDOUT.n63 VDDOUT.n56 416.101
R164 VDDOUT.n71 VDDOUT.n52 416.101
R165 VDDOUT.n74 VDDOUT.n48 416.101
R166 VDDOUT.n57 VDDOUT.n45 416.101
R167 VDDOUT.n42 VDDOUT.t3 356.894
R168 VDDOUT.n23 VDDOUT.n21 254.119
R169 VDDOUT.n37 VDDOUT.n4 254.119
R170 VDDOUT.n11 VDDOUT.n4 254.119
R171 VDDOUT.n12 VDDOUT.n11 254.119
R172 VDDOUT.n13 VDDOUT.n12 254.119
R173 VDDOUT.n7 VDDOUT.n1 254.119
R174 VDDOUT.n35 VDDOUT.n8 254.119
R175 VDDOUT.n31 VDDOUT.n8 254.119
R176 VDDOUT.n31 VDDOUT.n10 254.119
R177 VDDOUT.n27 VDDOUT.n10 254.119
R178 VDDOUT.n36 VDDOUT.n5 185.232
R179 VDDOUT.n28 VDDOUT.n14 185.232
R180 VDDOUT.n57 VDDOUT.n44 185
R181 VDDOUT.n57 VDDOUT.n55 185
R182 VDDOUT.n60 VDDOUT.n59 185
R183 VDDOUT.n61 VDDOUT.n56 185
R184 VDDOUT.n69 VDDOUT.n52 185
R185 VDDOUT.n52 VDDOUT.n51 185
R186 VDDOUT.n68 VDDOUT.n67 185
R187 VDDOUT.n67 VDDOUT.n66 185
R188 VDDOUT.n54 VDDOUT.n53 185
R189 VDDOUT.n65 VDDOUT.n54 185
R190 VDDOUT.n63 VDDOUT.n62 185
R191 VDDOUT.n64 VDDOUT.n63 185
R192 VDDOUT.n71 VDDOUT.n70 185
R193 VDDOUT.n50 VDDOUT.n49 185
R194 VDDOUT.n75 VDDOUT.n74 185
R195 VDDOUT.n74 VDDOUT.n73 185
R196 VDDOUT.n80 VDDOUT.n45 185
R197 VDDOUT.n64 VDDOUT.n45 185
R198 VDDOUT.n79 VDDOUT.n46 185
R199 VDDOUT.n65 VDDOUT.n46 185
R200 VDDOUT.n78 VDDOUT.n47 185
R201 VDDOUT.n66 VDDOUT.n47 185
R202 VDDOUT.n76 VDDOUT.n48 185
R203 VDDOUT.n51 VDDOUT.n48 185
R204 VDDOUT.n35 VDDOUT.n34 185
R205 VDDOUT.n36 VDDOUT.n35 185
R206 VDDOUT.n33 VDDOUT.n8 185
R207 VDDOUT.n8 VDDOUT.n6 185
R208 VDDOUT.n32 VDDOUT.n31 185
R209 VDDOUT.n31 VDDOUT.n30 185
R210 VDDOUT.n10 VDDOUT.n9 185
R211 VDDOUT.n29 VDDOUT.n10 185
R212 VDDOUT.n27 VDDOUT.n26 185
R213 VDDOUT.n28 VDDOUT.n27 185
R214 VDDOUT.n25 VDDOUT.n15 185
R215 VDDOUT.n24 VDDOUT.n23 185
R216 VDDOUT.n21 VDDOUT.n20 185
R217 VDDOUT.n21 VDDOUT.n14 185
R218 VDDOUT.n19 VDDOUT.n13 185
R219 VDDOUT.n28 VDDOUT.n13 185
R220 VDDOUT.n18 VDDOUT.n12 185
R221 VDDOUT.n29 VDDOUT.n12 185
R222 VDDOUT.n17 VDDOUT.n11 185
R223 VDDOUT.n30 VDDOUT.n11 185
R224 VDDOUT.n16 VDDOUT.n4 185
R225 VDDOUT.n6 VDDOUT.n4 185
R226 VDDOUT.n37 VDDOUT.n2 185
R227 VDDOUT.n37 VDDOUT.n36 185
R228 VDDOUT.n39 VDDOUT.n38 185
R229 VDDOUT.n40 VDDOUT.n1 185
R230 VDDOUT.n7 VDDOUT.n0 185
R231 VDDOUT.n7 VDDOUT.n5 185
R232 VDDOUT.n64 VDDOUT.n55 177.941
R233 VDDOUT.n73 VDDOUT.n51 177.941
R234 VDDOUT.n63 VDDOUT.n54 136.8
R235 VDDOUT.n67 VDDOUT.n54 136.8
R236 VDDOUT.n67 VDDOUT.n52 136.8
R237 VDDOUT.n74 VDDOUT.n50 136.8
R238 VDDOUT.n46 VDDOUT.n45 136.8
R239 VDDOUT.n47 VDDOUT.n46 136.8
R240 VDDOUT.n48 VDDOUT.n47 136.8
R241 VDDOUT.n59 VDDOUT.n57 136.8
R242 VDDOUT.n36 VDDOUT.n6 132.047
R243 VDDOUT.n30 VDDOUT.n29 132.047
R244 VDDOUT.n29 VDDOUT.n28 132.047
R245 VDDOUT.n65 VDDOUT.n64 105.882
R246 VDDOUT.n66 VDDOUT.n51 105.882
R247 VDDOUT.n22 VDDOUT.n15 75.3262
R248 VDDOUT.n38 VDDOUT.n3 75.3262
R249 VDDOUT.n23 VDDOUT.n22 75.3262
R250 VDDOUT.n3 VDDOUT.n1 75.3262
R251 VDDOUT.n26 VDDOUT.n25 72.6593
R252 VDDOUT.n20 VDDOUT.n19 72.6593
R253 VDDOUT.n39 VDDOUT.n2 72.6593
R254 VDDOUT.n34 VDDOUT.n0 72.2398
R255 VDDOUT.t2 VDDOUT.n6 69.6916
R256 VDDOUT.n58 VDDOUT.n55 67.5326
R257 VDDOUT.n73 VDDOUT.n72 67.5326
R258 VDDOUT.n30 VDDOUT.t2 62.3557
R259 VDDOUT.n22 VDDOUT.n14 54.8384
R260 VDDOUT.n5 VDDOUT.n3 54.8384
R261 VDDOUT.t0 VDDOUT.n65 52.9417
R262 VDDOUT.n66 VDDOUT.t0 52.9417
R263 VDDOUT.n72 VDDOUT.n71 49.9379
R264 VDDOUT.n59 VDDOUT.n58 49.9379
R265 VDDOUT.n58 VDDOUT.n56 49.9379
R266 VDDOUT.n72 VDDOUT.n50 49.9379
R267 VDDOUT.n80 VDDOUT.n44 46.7205
R268 VDDOUT.n62 VDDOUT.n61 46.7205
R269 VDDOUT.n70 VDDOUT.n69 46.7205
R270 VDDOUT.n76 VDDOUT.n75 46.7205
R271 VDDOUT.n34 VDDOUT.n33 27.1064
R272 VDDOUT.n33 VDDOUT.n32 27.1064
R273 VDDOUT.n32 VDDOUT.n9 27.1064
R274 VDDOUT.n26 VDDOUT.n9 27.1064
R275 VDDOUT.n25 VDDOUT.n24 27.1064
R276 VDDOUT.n24 VDDOUT.n20 27.1064
R277 VDDOUT.n16 VDDOUT.n2 27.1064
R278 VDDOUT.n17 VDDOUT.n16 27.1064
R279 VDDOUT.n18 VDDOUT.n17 27.1064
R280 VDDOUT.n19 VDDOUT.n18 27.1064
R281 VDDOUT.n40 VDDOUT.n39 26.6223
R282 VDDOUT.n60 VDDOUT.n44 15.3605
R283 VDDOUT.n61 VDDOUT.n60 15.3605
R284 VDDOUT.n62 VDDOUT.n53 15.3605
R285 VDDOUT.n68 VDDOUT.n53 15.3605
R286 VDDOUT.n69 VDDOUT.n68 15.3605
R287 VDDOUT.n75 VDDOUT.n49 15.3605
R288 VDDOUT.n70 VDDOUT.n49 15.3605
R289 VDDOUT.n80 VDDOUT.n79 15.3605
R290 VDDOUT.n79 VDDOUT.n78 15.3605
R291 VDDOUT.n81 VDDOUT.n80 9.3005
R292 VDDOUT.n79 VDDOUT.n43 9.3005
R293 VDDOUT.n41 VDDOUT.n40 5.52061
R294 VDDOUT.n41 VDDOUT.n0 5.433
R295 VDDOUT.n77 VDDOUT.n76 4.25641
R296 VDDOUT.n78 VDDOUT.n77 4.18886
R297 VDDOUT.n77 VDDOUT.n43 2.72752
R298 VDDOUT.n42 VDDOUT.n41 2.52943
R299 VDDOUT.n83 VDDOUT.n82 0.658833
R300 VDDOUT.n82 VDDOUT.n81 0.390083
R301 VDDOUT VDDOUT.n83 0.3385
R302 VDDOUT.n81 VDDOUT.n43 0.1505
R303 VDDOUT.n83 VDDOUT.n42 0.098
C0 IN VDDOUT 0.462527f
C1 IN a_259_346# 0.297618f
C2 IN OUT 0.011305f
C3 VDDOUT a_259_346# 0.623998f
C4 OUT VDDOUT 0.384118f
C5 OUT a_259_346# 0.246839f
C6 OUT VGND 0.59729f
C7 IN VGND 0.939247f
C8 VDDOUT VGND 4.48499f
C9 a_259_346# VGND 0.920816f
.ends

