** sch_path: /home/leo/Projects/IPs/sky130_leo_ip__levelshifter/xschem/sky130_leo_ip__levelshifter_up.sch
.subckt sky130_leo_ip__levelshifter_up VDDOUT VDDIN OUT IN VGND
*.PININFO IN:I VGND:B VDDIN:B OUT:I VDDOUT:B
XM1 ctrl_n IN VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 ctrl_n IN VDDIN VDDIN sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 ctrl ctrl_n VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 ctrl ctrl_n VDDIN VDDIN sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 OUT p1 VDDOUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM6 p1 ctrl VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 p1 OUT VDDOUT VDDOUT sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM8 OUT ctrl_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends
.end
