* NGSPICE file created from sky130_leo_ip__levelshifter_up.ext - technology: sky130A

.subckt sky130_leo_ip__levelshifter_up VDDOUT VDDIN OUT IN VGND
X0 VDDIN.t3 a_373_442# a_897_442# VDDIN.t2 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1 OUT.t1 a_373_442# VGND.t7 VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X2 VDDIN.t1 IN.t0 a_373_442# VDDIN.t0 sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X3 a_897_442# a_373_442# VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X4 VDDOUT.t3 OUT.t2 a_1778_346# VDDOUT.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X5 a_1778_346# a_897_442# VGND.t1 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X6 VDDOUT.t1 a_1778_346# OUT.t0 VDDOUT.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.5
X7 a_373_442# IN.t1 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
R0 VDDIN.n0 VDDIN.t2 473.38
R1 VDDIN.n1 VDDIN.n0 379.356
R2 VDDIN.n0 VDDIN.t0 376.11
R3 VDDIN.n2 VDDIN.t3 356.716
R4 VDDIN.n1 VDDIN.t1 356.635
R5 VDDIN VDDIN.n2 0.3385
R6 VDDIN.n2 VDDIN.n1 0.00425
R7 VGND.n329 VGND.n328 5095.62
R8 VGND.n331 VGND.n54 1980
R9 VGND.n339 VGND.n54 1980
R10 VGND.n340 VGND.n339 1980
R11 VGND.n341 VGND.n340 1980
R12 VGND.n341 VGND.n48 1980
R13 VGND.n349 VGND.n48 1980
R14 VGND.n350 VGND.n349 1980
R15 VGND.n351 VGND.n350 1980
R16 VGND.n351 VGND.n41 1980
R17 VGND.n361 VGND.n41 1980
R18 VGND.n362 VGND.n361 1980
R19 VGND.n363 VGND.n362 1980
R20 VGND.n38 VGND.n33 1766.93
R21 VGND.n374 VGND.n33 1247.24
R22 VGND.n375 VGND.n374 1247.24
R23 VGND.n376 VGND.n375 1247.24
R24 VGND.n376 VGND.n27 1247.24
R25 VGND.n384 VGND.n27 1247.24
R26 VGND.n385 VGND.n384 1247.24
R27 VGND.n386 VGND.n385 1247.24
R28 VGND.n133 VGND.n131 1152
R29 VGND.n134 VGND.n133 1152
R30 VGND.n135 VGND.n134 1152
R31 VGND.n136 VGND.n135 1152
R32 VGND.n138 VGND.n136 1152
R33 VGND.n139 VGND.n138 1152
R34 VGND.n140 VGND.n139 1152
R35 VGND.n141 VGND.n140 1152
R36 VGND.n142 VGND.n141 1152
R37 VGND.n143 VGND.n142 1152
R38 VGND.n143 VGND.n61 1152
R39 VGND.n114 VGND.n109 1112.5
R40 VGND.n331 VGND.n330 1100
R41 VGND.n363 VGND.n38 1100
R42 VGND.n386 VGND.n16 1039.37
R43 VGND.n193 VGND.n192 900
R44 VGND.n194 VGND.n193 900
R45 VGND.n194 VGND.n103 900
R46 VGND.n202 VGND.n103 900
R47 VGND.n203 VGND.n202 900
R48 VGND.n204 VGND.n203 900
R49 VGND.n204 VGND.n95 900
R50 VGND.n231 VGND.n95 900
R51 VGND.n232 VGND.n231 837.5
R52 VGND.n367 VGND.n34 800.848
R53 VGND.n407 VGND.n13 800.848
R54 VGND.n234 VGND.n93 800.848
R55 VGND.n191 VGND.n110 800.848
R56 VGND.n366 VGND.n38 768.5
R57 VGND.n111 VGND.n110 585
R58 VGND.n114 VGND.n110 585
R59 VGND.n186 VGND.n113 585
R60 VGND.n185 VGND.n116 585
R61 VGND.n184 VGND.n117 585
R62 VGND.n131 VGND.n117 585
R63 VGND.n132 VGND.n118 585
R64 VGND.n133 VGND.n132 585
R65 VGND.n180 VGND.n120 585
R66 VGND.n134 VGND.n120 585
R67 VGND.n179 VGND.n121 585
R68 VGND.n135 VGND.n121 585
R69 VGND.n178 VGND.n122 585
R70 VGND.n136 VGND.n122 585
R71 VGND.n137 VGND.n123 585
R72 VGND.n138 VGND.n137 585
R73 VGND.n174 VGND.n125 585
R74 VGND.n139 VGND.n125 585
R75 VGND.n173 VGND.n126 585
R76 VGND.n140 VGND.n126 585
R77 VGND.n172 VGND.n127 585
R78 VGND.n141 VGND.n127 585
R79 VGND.n130 VGND.n128 585
R80 VGND.n142 VGND.n130 585
R81 VGND.n168 VGND.n144 585
R82 VGND.n144 VGND.n143 585
R83 VGND.n167 VGND.n145 585
R84 VGND.n145 VGND.n61 585
R85 VGND.n166 VGND.n146 585
R86 VGND.n150 VGND.n147 585
R87 VGND.n162 VGND.n151 585
R88 VGND.n161 VGND.n153 585
R89 VGND.n160 VGND.n154 585
R90 VGND.n157 VGND.n156 585
R91 VGND.n59 VGND.n58 585
R92 VGND.n60 VGND.n59 585
R93 VGND.n333 VGND.n332 585
R94 VGND.n332 VGND.n331 585
R95 VGND.n56 VGND.n55 585
R96 VGND.n55 VGND.n54 585
R97 VGND.n338 VGND.n337 585
R98 VGND.n339 VGND.n338 585
R99 VGND.n53 VGND.n52 585
R100 VGND.n340 VGND.n53 585
R101 VGND.n343 VGND.n342 585
R102 VGND.n342 VGND.n341 585
R103 VGND.n50 VGND.n49 585
R104 VGND.n49 VGND.n48 585
R105 VGND.n348 VGND.n347 585
R106 VGND.n349 VGND.n348 585
R107 VGND.n47 VGND.n46 585
R108 VGND.n350 VGND.n47 585
R109 VGND.n353 VGND.n352 585
R110 VGND.n352 VGND.n351 585
R111 VGND.n43 VGND.n42 585
R112 VGND.n42 VGND.n41 585
R113 VGND.n360 VGND.n359 585
R114 VGND.n361 VGND.n360 585
R115 VGND.n44 VGND.n39 585
R116 VGND.n362 VGND.n39 585
R117 VGND.n364 VGND.n40 585
R118 VGND.n364 VGND.n363 585
R119 VGND.n365 VGND.n37 585
R120 VGND.n368 VGND.n367 585
R121 VGND.n191 VGND.n190 585
R122 VGND.n192 VGND.n191 585
R123 VGND.n108 VGND.n107 585
R124 VGND.n193 VGND.n108 585
R125 VGND.n196 VGND.n195 585
R126 VGND.n195 VGND.n194 585
R127 VGND.n105 VGND.n104 585
R128 VGND.n104 VGND.n103 585
R129 VGND.n201 VGND.n200 585
R130 VGND.n202 VGND.n201 585
R131 VGND.n102 VGND.n101 585
R132 VGND.n203 VGND.n102 585
R133 VGND.n206 VGND.n205 585
R134 VGND.n205 VGND.n204 585
R135 VGND.n98 VGND.n96 585
R136 VGND.n96 VGND.n95 585
R137 VGND.n230 VGND.n229 585
R138 VGND.n231 VGND.n230 585
R139 VGND.n99 VGND.n97 585
R140 VGND.n225 VGND.n211 585
R141 VGND.n224 VGND.n212 585
R142 VGND.n212 VGND.n94 585
R143 VGND.n223 VGND.n213 585
R144 VGND.n216 VGND.n214 585
R145 VGND.n219 VGND.n218 585
R146 VGND.n93 VGND.n92 585
R147 VGND.n409 VGND.n13 585
R148 VGND.n296 VGND.n13 585
R149 VGND.n297 VGND.n11 585
R150 VGND.n298 VGND.n297 585
R151 VGND.n413 VGND.n10 585
R152 VGND.n299 VGND.n10 585
R153 VGND.n414 VGND.n9 585
R154 VGND.n300 VGND.n9 585
R155 VGND.n415 VGND.n8 585
R156 VGND.n301 VGND.n8 585
R157 VGND.n302 VGND.n6 585
R158 VGND.n303 VGND.n302 585
R159 VGND.n420 VGND.n5 585
R160 VGND.n304 VGND.n5 585
R161 VGND.n421 VGND.n4 585
R162 VGND.n305 VGND.n4 585
R163 VGND.n422 VGND.n3 585
R164 VGND.n306 VGND.n3 585
R165 VGND.n288 VGND.n2 585
R166 VGND.n307 VGND.n288 585
R167 VGND.n310 VGND.n309 585
R168 VGND.n309 VGND.n308 585
R169 VGND.n313 VGND.n287 585
R170 VGND.n295 VGND.n287 585
R171 VGND.n314 VGND.n286 585
R172 VGND.n294 VGND.n286 585
R173 VGND.n292 VGND.n284 585
R174 VGND.n293 VGND.n292 585
R175 VGND.n318 VGND.n283 585
R176 VGND.n291 VGND.n283 585
R177 VGND.n319 VGND.n282 585
R178 VGND.n290 VGND.n282 585
R179 VGND.n320 VGND.n281 585
R180 VGND.n289 VGND.n281 585
R181 VGND.n67 VGND.n65 585
R182 VGND.n65 VGND.n63 585
R183 VGND.n326 VGND.n325 585
R184 VGND.n327 VGND.n326 585
R185 VGND.n66 VGND.n64 585
R186 VGND.n64 VGND.n62 585
R187 VGND.n276 VGND.n275 585
R188 VGND.n275 VGND.n274 585
R189 VGND.n70 VGND.n69 585
R190 VGND.n273 VGND.n70 585
R191 VGND.n271 VGND.n270 585
R192 VGND.n272 VGND.n271 585
R193 VGND.n73 VGND.n72 585
R194 VGND.n72 VGND.n71 585
R195 VGND.n266 VGND.n265 585
R196 VGND.n265 VGND.n264 585
R197 VGND.n76 VGND.n75 585
R198 VGND.n263 VGND.n76 585
R199 VGND.n261 VGND.n260 585
R200 VGND.n262 VGND.n261 585
R201 VGND.n79 VGND.n78 585
R202 VGND.n78 VGND.n77 585
R203 VGND.n256 VGND.n255 585
R204 VGND.n255 VGND.n254 585
R205 VGND.n82 VGND.n81 585
R206 VGND.n253 VGND.n82 585
R207 VGND.n251 VGND.n250 585
R208 VGND.n252 VGND.n251 585
R209 VGND.n84 VGND.n83 585
R210 VGND.n243 VGND.n83 585
R211 VGND.n246 VGND.n245 585
R212 VGND.n245 VGND.n244 585
R213 VGND.n87 VGND.n86 585
R214 VGND.n242 VGND.n87 585
R215 VGND.n240 VGND.n239 585
R216 VGND.n241 VGND.n240 585
R217 VGND.n90 VGND.n89 585
R218 VGND.n89 VGND.n88 585
R219 VGND.n235 VGND.n234 585
R220 VGND.n234 VGND.n233 585
R221 VGND.n408 VGND.n407 585
R222 VGND.n15 VGND.n14 585
R223 VGND.n403 VGND.n402 585
R224 VGND.n20 VGND.n19 585
R225 VGND.n397 VGND.n396 585
R226 VGND.n395 VGND.n394 585
R227 VGND.n393 VGND.n392 585
R228 VGND.n26 VGND.n22 585
R229 VGND.n388 VGND.n387 585
R230 VGND.n387 VGND.n386 585
R231 VGND.n25 VGND.n24 585
R232 VGND.n385 VGND.n25 585
R233 VGND.n383 VGND.n382 585
R234 VGND.n384 VGND.n383 585
R235 VGND.n29 VGND.n28 585
R236 VGND.n28 VGND.n27 585
R237 VGND.n378 VGND.n377 585
R238 VGND.n377 VGND.n376 585
R239 VGND.n32 VGND.n31 585
R240 VGND.n375 VGND.n32 585
R241 VGND.n373 VGND.n372 585
R242 VGND.n374 VGND.n373 585
R243 VGND.n35 VGND.n34 585
R244 VGND.n34 VGND.n33 585
R245 VGND.n192 VGND.n109 550
R246 VGND.n233 VGND.n94 547.335
R247 VGND.n241 VGND.n88 511.793
R248 VGND.n242 VGND.n241 511.793
R249 VGND.n244 VGND.n242 511.793
R250 VGND.n244 VGND.n243 511.793
R251 VGND.n253 VGND.n252 511.793
R252 VGND.n254 VGND.n253 511.793
R253 VGND.n254 VGND.n77 511.793
R254 VGND.n262 VGND.n77 511.793
R255 VGND.n263 VGND.n262 511.793
R256 VGND.n264 VGND.n71 511.793
R257 VGND.n272 VGND.n71 511.793
R258 VGND.n330 VGND.n329 486.096
R259 VGND.n273 VGND.n272 462.719
R260 VGND.n274 VGND.n273 453.868
R261 VGND.n274 VGND.n62 453.868
R262 VGND.n327 VGND.n63 453.868
R263 VGND.n289 VGND.n63 453.868
R264 VGND.n290 VGND.n289 453.868
R265 VGND.n291 VGND.n290 453.868
R266 VGND.n293 VGND.n291 453.868
R267 VGND.n294 VGND.n293 453.868
R268 VGND.n308 VGND.n295 453.868
R269 VGND.n308 VGND.n307 453.868
R270 VGND.n307 VGND.n306 453.868
R271 VGND.n306 VGND.n305 453.868
R272 VGND.n305 VGND.n304 453.868
R273 VGND.n304 VGND.n303 453.868
R274 VGND.n301 VGND.n300 453.868
R275 VGND.n300 VGND.n299 453.868
R276 VGND.n299 VGND.n298 453.868
R277 VGND.n298 VGND.n296 453.868
R278 VGND.n303 VGND.t2 441.262
R279 VGND.n232 VGND.n88 405.171
R280 VGND.n243 VGND.t6 405.171
R281 VGND.n131 VGND.n109 400
R282 VGND.n328 VGND.n62 365.616
R283 VGND.n405 VGND.n16 340.401
R284 VGND.t0 VGND.n263 334.087
R285 VGND.t4 VGND.n294 315.187
R286 VGND.n373 VGND.n34 308.349
R287 VGND.n373 VGND.n32 308.349
R288 VGND.n377 VGND.n32 308.349
R289 VGND.n377 VGND.n28 308.349
R290 VGND.n383 VGND.n28 308.349
R291 VGND.n383 VGND.n25 308.349
R292 VGND.n387 VGND.n25 308.349
R293 VGND.n387 VGND.n26 308.349
R294 VGND.n394 VGND.n393 308.349
R295 VGND.n396 VGND.n19 308.349
R296 VGND.n403 VGND.n15 308.349
R297 VGND.n234 VGND.n89 308.349
R298 VGND.n240 VGND.n89 308.349
R299 VGND.n240 VGND.n87 308.349
R300 VGND.n245 VGND.n87 308.349
R301 VGND.n245 VGND.n83 308.349
R302 VGND.n251 VGND.n83 308.349
R303 VGND.n251 VGND.n82 308.349
R304 VGND.n255 VGND.n82 308.349
R305 VGND.n255 VGND.n78 308.349
R306 VGND.n261 VGND.n78 308.349
R307 VGND.n261 VGND.n76 308.349
R308 VGND.n265 VGND.n76 308.349
R309 VGND.n265 VGND.n72 308.349
R310 VGND.n271 VGND.n72 308.349
R311 VGND.n271 VGND.n70 308.349
R312 VGND.n275 VGND.n70 308.349
R313 VGND.n275 VGND.n64 308.349
R314 VGND.n326 VGND.n64 308.349
R315 VGND.n326 VGND.n65 308.349
R316 VGND.n281 VGND.n65 308.349
R317 VGND.n282 VGND.n281 308.349
R318 VGND.n283 VGND.n282 308.349
R319 VGND.n292 VGND.n283 308.349
R320 VGND.n292 VGND.n286 308.349
R321 VGND.n287 VGND.n286 308.349
R322 VGND.n309 VGND.n287 308.349
R323 VGND.n309 VGND.n288 308.349
R324 VGND.n288 VGND.n3 308.349
R325 VGND.n4 VGND.n3 308.349
R326 VGND.n5 VGND.n4 308.349
R327 VGND.n302 VGND.n5 308.349
R328 VGND.n302 VGND.n8 308.349
R329 VGND.n9 VGND.n8 308.349
R330 VGND.n10 VGND.n9 308.349
R331 VGND.n297 VGND.n10 308.349
R332 VGND.n297 VGND.n13 308.349
R333 VGND.n191 VGND.n108 308.349
R334 VGND.n195 VGND.n108 308.349
R335 VGND.n195 VGND.n104 308.349
R336 VGND.n201 VGND.n104 308.349
R337 VGND.n201 VGND.n102 308.349
R338 VGND.n205 VGND.n102 308.349
R339 VGND.n205 VGND.n96 308.349
R340 VGND.n230 VGND.n96 308.349
R341 VGND.n230 VGND.n97 308.349
R342 VGND.n212 VGND.n211 308.349
R343 VGND.n213 VGND.n212 308.349
R344 VGND.n218 VGND.n216 308.349
R345 VGND.n113 VGND.n110 308.349
R346 VGND.n117 VGND.n116 308.349
R347 VGND.n132 VGND.n117 308.349
R348 VGND.n132 VGND.n120 308.349
R349 VGND.n121 VGND.n120 308.349
R350 VGND.n122 VGND.n121 308.349
R351 VGND.n137 VGND.n122 308.349
R352 VGND.n137 VGND.n125 308.349
R353 VGND.n126 VGND.n125 308.349
R354 VGND.n127 VGND.n126 308.349
R355 VGND.n130 VGND.n127 308.349
R356 VGND.n144 VGND.n130 308.349
R357 VGND.n145 VGND.n144 308.349
R358 VGND.n146 VGND.n145 308.349
R359 VGND.n151 VGND.n150 308.349
R360 VGND.n154 VGND.n153 308.349
R361 VGND.n156 VGND.n59 308.349
R362 VGND.n332 VGND.n59 308.349
R363 VGND.n332 VGND.n55 308.349
R364 VGND.n338 VGND.n55 308.349
R365 VGND.n338 VGND.n53 308.349
R366 VGND.n342 VGND.n53 308.349
R367 VGND.n342 VGND.n49 308.349
R368 VGND.n348 VGND.n49 308.349
R369 VGND.n348 VGND.n47 308.349
R370 VGND.n352 VGND.n47 308.349
R371 VGND.n352 VGND.n42 308.349
R372 VGND.n360 VGND.n42 308.349
R373 VGND.n360 VGND.n39 308.349
R374 VGND.n364 VGND.n39 308.349
R375 VGND.n365 VGND.n364 308.349
R376 VGND.n330 VGND.n60 259.81
R377 VGND.n285 VGND.t5 237.345
R378 VGND.n417 VGND.t3 237.345
R379 VGND.n115 VGND.n114 231.493
R380 VGND.n149 VGND.n60 231.493
R381 VGND.n152 VGND.n60 231.493
R382 VGND.n155 VGND.n60 231.493
R383 VGND.n210 VGND.n94 231.493
R384 VGND.n215 VGND.n94 231.493
R385 VGND.n217 VGND.n94 231.493
R386 VGND.n406 VGND.n405 231.493
R387 VGND.n405 VGND.n404 231.493
R388 VGND.n405 VGND.n18 231.493
R389 VGND.n405 VGND.n17 231.493
R390 VGND.n264 VGND.t0 177.707
R391 VGND.n329 VGND.n61 176
R392 VGND.n296 VGND.n16 144.987
R393 VGND.n295 VGND.t4 138.683
R394 VGND.n279 VGND.t7 131.897
R395 VGND.n279 VGND.t1 131.332
R396 VGND.n393 VGND.n17 122.017
R397 VGND.n396 VGND.n18 122.017
R398 VGND.n404 VGND.n403 122.017
R399 VGND.n407 VGND.n406 122.017
R400 VGND.n210 VGND.n97 122.017
R401 VGND.n215 VGND.n213 122.017
R402 VGND.n218 VGND.n217 122.017
R403 VGND.n116 VGND.n115 122.017
R404 VGND.n149 VGND.n146 122.017
R405 VGND.n152 VGND.n151 122.017
R406 VGND.n155 VGND.n154 122.017
R407 VGND.n366 VGND.n365 122.017
R408 VGND.n115 VGND.n113 122.017
R409 VGND.n150 VGND.n149 122.017
R410 VGND.n153 VGND.n152 122.017
R411 VGND.n156 VGND.n155 122.017
R412 VGND.n367 VGND.n366 122.017
R413 VGND.n211 VGND.n210 122.017
R414 VGND.n216 VGND.n215 122.017
R415 VGND.n217 VGND.n93 122.017
R416 VGND.n406 VGND.n15 122.017
R417 VGND.n404 VGND.n19 122.017
R418 VGND.n394 VGND.n18 122.017
R419 VGND.n26 VGND.n17 122.017
R420 VGND.n233 VGND.n232 106.624
R421 VGND.n252 VGND.t6 106.624
R422 VGND.n328 VGND.n327 88.2527
R423 VGND.n190 VGND.n111 52.0353
R424 VGND.n368 VGND.n35 52.0353
R425 VGND.n235 VGND.n92 52.0353
R426 VGND.n409 VGND.n408 52.0353
R427 VGND.n186 VGND.n111 20.0353
R428 VGND.n186 VGND.n185 20.0353
R429 VGND.n185 VGND.n184 20.0353
R430 VGND.n184 VGND.n118 20.0353
R431 VGND.n180 VGND.n118 20.0353
R432 VGND.n180 VGND.n179 20.0353
R433 VGND.n179 VGND.n178 20.0353
R434 VGND.n178 VGND.n123 20.0353
R435 VGND.n174 VGND.n123 20.0353
R436 VGND.n174 VGND.n173 20.0353
R437 VGND.n173 VGND.n172 20.0353
R438 VGND.n172 VGND.n128 20.0353
R439 VGND.n168 VGND.n128 20.0353
R440 VGND.n168 VGND.n167 20.0353
R441 VGND.n167 VGND.n166 20.0353
R442 VGND.n166 VGND.n147 20.0353
R443 VGND.n162 VGND.n147 20.0353
R444 VGND.n162 VGND.n161 20.0353
R445 VGND.n161 VGND.n160 20.0353
R446 VGND.n160 VGND.n157 20.0353
R447 VGND.n157 VGND.n58 20.0353
R448 VGND.n333 VGND.n58 20.0353
R449 VGND.n333 VGND.n56 20.0353
R450 VGND.n337 VGND.n56 20.0353
R451 VGND.n337 VGND.n52 20.0353
R452 VGND.n343 VGND.n52 20.0353
R453 VGND.n343 VGND.n50 20.0353
R454 VGND.n347 VGND.n50 20.0353
R455 VGND.n347 VGND.n46 20.0353
R456 VGND.n353 VGND.n46 20.0353
R457 VGND.n353 VGND.n43 20.0353
R458 VGND.n359 VGND.n43 20.0353
R459 VGND.n359 VGND.n44 20.0353
R460 VGND.n44 VGND.n40 20.0353
R461 VGND.n40 VGND.n37 20.0353
R462 VGND.n368 VGND.n37 20.0353
R463 VGND.n190 VGND.n107 20.0353
R464 VGND.n196 VGND.n107 20.0353
R465 VGND.n196 VGND.n105 20.0353
R466 VGND.n200 VGND.n105 20.0353
R467 VGND.n200 VGND.n101 20.0353
R468 VGND.n206 VGND.n101 20.0353
R469 VGND.n206 VGND.n98 20.0353
R470 VGND.n229 VGND.n98 20.0353
R471 VGND.n229 VGND.n99 20.0353
R472 VGND.n225 VGND.n99 20.0353
R473 VGND.n225 VGND.n224 20.0353
R474 VGND.n224 VGND.n223 20.0353
R475 VGND.n223 VGND.n214 20.0353
R476 VGND.n219 VGND.n214 20.0353
R477 VGND.n219 VGND.n92 20.0353
R478 VGND.n235 VGND.n90 20.0353
R479 VGND.n239 VGND.n90 20.0353
R480 VGND.n239 VGND.n86 20.0353
R481 VGND.n246 VGND.n86 20.0353
R482 VGND.n246 VGND.n84 20.0353
R483 VGND.n250 VGND.n84 20.0353
R484 VGND.n250 VGND.n81 20.0353
R485 VGND.n256 VGND.n81 20.0353
R486 VGND.n256 VGND.n79 20.0353
R487 VGND.n260 VGND.n79 20.0353
R488 VGND.n260 VGND.n75 20.0353
R489 VGND.n266 VGND.n75 20.0353
R490 VGND.n266 VGND.n73 20.0353
R491 VGND.n270 VGND.n73 20.0353
R492 VGND.n270 VGND.n69 20.0353
R493 VGND.n276 VGND.n69 20.0353
R494 VGND.n276 VGND.n66 20.0353
R495 VGND.n325 VGND.n66 20.0353
R496 VGND.n325 VGND.n67 20.0353
R497 VGND.n320 VGND.n67 20.0353
R498 VGND.n320 VGND.n319 20.0353
R499 VGND.n319 VGND.n318 20.0353
R500 VGND.n318 VGND.n284 20.0353
R501 VGND.n314 VGND.n284 20.0353
R502 VGND.n314 VGND.n313 20.0353
R503 VGND.n313 VGND.n310 20.0353
R504 VGND.n310 VGND.n2 20.0353
R505 VGND.n422 VGND.n2 20.0353
R506 VGND.n422 VGND.n421 20.0353
R507 VGND.n421 VGND.n420 20.0353
R508 VGND.n420 VGND.n6 20.0353
R509 VGND.n415 VGND.n6 20.0353
R510 VGND.n415 VGND.n414 20.0353
R511 VGND.n414 VGND.n413 20.0353
R512 VGND.n413 VGND.n11 20.0353
R513 VGND.n409 VGND.n11 20.0353
R514 VGND.n372 VGND.n35 20.0353
R515 VGND.n372 VGND.n31 20.0353
R516 VGND.n378 VGND.n31 20.0353
R517 VGND.n378 VGND.n29 20.0353
R518 VGND.n382 VGND.n29 20.0353
R519 VGND.n382 VGND.n24 20.0353
R520 VGND.n388 VGND.n24 20.0353
R521 VGND.n388 VGND.n22 20.0353
R522 VGND.n392 VGND.n22 20.0353
R523 VGND.n395 VGND.n392 20.0353
R524 VGND.n397 VGND.n395 20.0353
R525 VGND.n397 VGND.n20 20.0353
R526 VGND.n402 VGND.n20 20.0353
R527 VGND.n402 VGND.n14 20.0353
R528 VGND.n408 VGND.n14 20.0353
R529 VGND.t2 VGND.n301 12.608
R530 VGND.n408 VGND.n12 9.3005
R531 VGND.n400 VGND.n14 9.3005
R532 VGND.n402 VGND.n401 9.3005
R533 VGND.n399 VGND.n20 9.3005
R534 VGND.n398 VGND.n397 9.3005
R535 VGND.n395 VGND.n21 9.3005
R536 VGND.n392 VGND.n391 9.3005
R537 VGND.n390 VGND.n22 9.3005
R538 VGND.n389 VGND.n388 9.3005
R539 VGND.n24 VGND.n23 9.3005
R540 VGND.n382 VGND.n381 9.3005
R541 VGND.n380 VGND.n29 9.3005
R542 VGND.n379 VGND.n378 9.3005
R543 VGND.n31 VGND.n30 9.3005
R544 VGND.n372 VGND.n371 9.3005
R545 VGND.n370 VGND.n35 9.3005
R546 VGND.n188 VGND.n111 9.3005
R547 VGND.n187 VGND.n186 9.3005
R548 VGND.n185 VGND.n112 9.3005
R549 VGND.n184 VGND.n183 9.3005
R550 VGND.n182 VGND.n118 9.3005
R551 VGND.n181 VGND.n180 9.3005
R552 VGND.n179 VGND.n119 9.3005
R553 VGND.n178 VGND.n177 9.3005
R554 VGND.n176 VGND.n123 9.3005
R555 VGND.n175 VGND.n174 9.3005
R556 VGND.n173 VGND.n124 9.3005
R557 VGND.n172 VGND.n171 9.3005
R558 VGND.n170 VGND.n128 9.3005
R559 VGND.n169 VGND.n168 9.3005
R560 VGND.n167 VGND.n129 9.3005
R561 VGND.n166 VGND.n165 9.3005
R562 VGND.n164 VGND.n147 9.3005
R563 VGND.n163 VGND.n162 9.3005
R564 VGND.n161 VGND.n148 9.3005
R565 VGND.n160 VGND.n159 9.3005
R566 VGND.n158 VGND.n157 9.3005
R567 VGND.n58 VGND.n57 9.3005
R568 VGND.n334 VGND.n333 9.3005
R569 VGND.n335 VGND.n56 9.3005
R570 VGND.n337 VGND.n336 9.3005
R571 VGND.n52 VGND.n51 9.3005
R572 VGND.n344 VGND.n343 9.3005
R573 VGND.n345 VGND.n50 9.3005
R574 VGND.n347 VGND.n346 9.3005
R575 VGND.n46 VGND.n45 9.3005
R576 VGND.n354 VGND.n353 9.3005
R577 VGND.n355 VGND.n43 9.3005
R578 VGND.n359 VGND.n358 9.3005
R579 VGND.n357 VGND.n44 9.3005
R580 VGND.n356 VGND.n40 9.3005
R581 VGND.n37 VGND.n36 9.3005
R582 VGND.n369 VGND.n368 9.3005
R583 VGND.n190 VGND.n189 9.3005
R584 VGND.n107 VGND.n106 9.3005
R585 VGND.n197 VGND.n196 9.3005
R586 VGND.n198 VGND.n105 9.3005
R587 VGND.n200 VGND.n199 9.3005
R588 VGND.n101 VGND.n100 9.3005
R589 VGND.n207 VGND.n206 9.3005
R590 VGND.n208 VGND.n98 9.3005
R591 VGND.n229 VGND.n228 9.3005
R592 VGND.n227 VGND.n99 9.3005
R593 VGND.n226 VGND.n225 9.3005
R594 VGND.n224 VGND.n209 9.3005
R595 VGND.n223 VGND.n222 9.3005
R596 VGND.n221 VGND.n214 9.3005
R597 VGND.n220 VGND.n219 9.3005
R598 VGND.n92 VGND.n91 9.3005
R599 VGND.n323 VGND.n67 9.3005
R600 VGND.n325 VGND.n324 9.3005
R601 VGND.n278 VGND.n66 9.3005
R602 VGND.n277 VGND.n276 9.3005
R603 VGND.n69 VGND.n68 9.3005
R604 VGND.n270 VGND.n269 9.3005
R605 VGND.n268 VGND.n73 9.3005
R606 VGND.n267 VGND.n266 9.3005
R607 VGND.n75 VGND.n74 9.3005
R608 VGND.n260 VGND.n259 9.3005
R609 VGND.n258 VGND.n79 9.3005
R610 VGND.n257 VGND.n256 9.3005
R611 VGND.n81 VGND.n80 9.3005
R612 VGND.n250 VGND.n249 9.3005
R613 VGND.n248 VGND.n84 9.3005
R614 VGND.n247 VGND.n246 9.3005
R615 VGND.n86 VGND.n85 9.3005
R616 VGND.n239 VGND.n238 9.3005
R617 VGND.n237 VGND.n90 9.3005
R618 VGND.n236 VGND.n235 9.3005
R619 VGND.n410 VGND.n409 9.3005
R620 VGND.n411 VGND.n11 9.3005
R621 VGND.n413 VGND.n412 9.3005
R622 VGND.n414 VGND.n7 9.3005
R623 VGND.n416 VGND.n415 9.3005
R624 VGND.n418 VGND.n6 9.3005
R625 VGND.n420 VGND.n419 9.3005
R626 VGND.n421 VGND.n1 9.3005
R627 VGND.n423 VGND.n422 9.3005
R628 VGND.n2 VGND.n0 9.3005
R629 VGND.n311 VGND.n310 9.3005
R630 VGND.n313 VGND.n312 9.3005
R631 VGND.n315 VGND.n314 9.3005
R632 VGND.n316 VGND.n284 9.3005
R633 VGND.n318 VGND.n317 9.3005
R634 VGND.n319 VGND.n280 9.3005
R635 VGND.n321 VGND.n320 9.3005
R636 VGND.n322 VGND.n279 0.798406
R637 VGND.n370 VGND.n369 0.508652
R638 VGND.n189 VGND.n188 0.508652
R639 VGND.n236 VGND.n91 0.508652
R640 VGND.n410 VGND.n12 0.470327
R641 VGND VGND.n424 0.3385
R642 VGND.n371 VGND.n370 0.196152
R643 VGND.n371 VGND.n30 0.196152
R644 VGND.n379 VGND.n30 0.196152
R645 VGND.n380 VGND.n379 0.196152
R646 VGND.n381 VGND.n380 0.196152
R647 VGND.n381 VGND.n23 0.196152
R648 VGND.n389 VGND.n23 0.196152
R649 VGND.n390 VGND.n389 0.196152
R650 VGND.n391 VGND.n390 0.196152
R651 VGND.n391 VGND.n21 0.196152
R652 VGND.n398 VGND.n21 0.196152
R653 VGND.n399 VGND.n398 0.196152
R654 VGND.n401 VGND.n399 0.196152
R655 VGND.n401 VGND.n400 0.196152
R656 VGND.n400 VGND.n12 0.196152
R657 VGND.n188 VGND.n187 0.196152
R658 VGND.n187 VGND.n112 0.196152
R659 VGND.n183 VGND.n112 0.196152
R660 VGND.n183 VGND.n182 0.196152
R661 VGND.n182 VGND.n181 0.196152
R662 VGND.n181 VGND.n119 0.196152
R663 VGND.n177 VGND.n119 0.196152
R664 VGND.n177 VGND.n176 0.196152
R665 VGND.n176 VGND.n175 0.196152
R666 VGND.n175 VGND.n124 0.196152
R667 VGND.n171 VGND.n124 0.196152
R668 VGND.n171 VGND.n170 0.196152
R669 VGND.n170 VGND.n169 0.196152
R670 VGND.n169 VGND.n129 0.196152
R671 VGND.n165 VGND.n129 0.196152
R672 VGND.n165 VGND.n164 0.196152
R673 VGND.n164 VGND.n163 0.196152
R674 VGND.n163 VGND.n148 0.196152
R675 VGND.n159 VGND.n148 0.196152
R676 VGND.n159 VGND.n158 0.196152
R677 VGND.n158 VGND.n57 0.196152
R678 VGND.n334 VGND.n57 0.196152
R679 VGND.n335 VGND.n334 0.196152
R680 VGND.n336 VGND.n335 0.196152
R681 VGND.n336 VGND.n51 0.196152
R682 VGND.n344 VGND.n51 0.196152
R683 VGND.n345 VGND.n344 0.196152
R684 VGND.n346 VGND.n345 0.196152
R685 VGND.n346 VGND.n45 0.196152
R686 VGND.n354 VGND.n45 0.196152
R687 VGND.n355 VGND.n354 0.196152
R688 VGND.n358 VGND.n355 0.196152
R689 VGND.n358 VGND.n357 0.196152
R690 VGND.n357 VGND.n356 0.196152
R691 VGND.n356 VGND.n36 0.196152
R692 VGND.n369 VGND.n36 0.196152
R693 VGND.n189 VGND.n106 0.196152
R694 VGND.n197 VGND.n106 0.196152
R695 VGND.n198 VGND.n197 0.196152
R696 VGND.n199 VGND.n198 0.196152
R697 VGND.n199 VGND.n100 0.196152
R698 VGND.n207 VGND.n100 0.196152
R699 VGND.n208 VGND.n207 0.196152
R700 VGND.n228 VGND.n208 0.196152
R701 VGND.n228 VGND.n227 0.196152
R702 VGND.n227 VGND.n226 0.196152
R703 VGND.n226 VGND.n209 0.196152
R704 VGND.n222 VGND.n209 0.196152
R705 VGND.n222 VGND.n221 0.196152
R706 VGND.n221 VGND.n220 0.196152
R707 VGND.n220 VGND.n91 0.196152
R708 VGND.n237 VGND.n236 0.196152
R709 VGND.n238 VGND.n237 0.196152
R710 VGND.n238 VGND.n85 0.196152
R711 VGND.n247 VGND.n85 0.196152
R712 VGND.n248 VGND.n247 0.196152
R713 VGND.n249 VGND.n248 0.196152
R714 VGND.n249 VGND.n80 0.196152
R715 VGND.n257 VGND.n80 0.196152
R716 VGND.n258 VGND.n257 0.196152
R717 VGND.n259 VGND.n258 0.196152
R718 VGND.n259 VGND.n74 0.196152
R719 VGND.n267 VGND.n74 0.196152
R720 VGND.n268 VGND.n267 0.196152
R721 VGND.n269 VGND.n268 0.196152
R722 VGND.n269 VGND.n68 0.196152
R723 VGND.n277 VGND.n68 0.196152
R724 VGND.n278 VGND.n277 0.196152
R725 VGND.n324 VGND.n278 0.196152
R726 VGND.n324 VGND.n323 0.196152
R727 VGND.n323 VGND.n322 0.111913
R728 VGND.n321 VGND.n280 0.0338333
R729 VGND.n317 VGND.n280 0.0338333
R730 VGND.n317 VGND.n316 0.0338333
R731 VGND.n316 VGND.n315 0.0338333
R732 VGND.n312 VGND.n311 0.0338333
R733 VGND.n311 VGND.n0 0.0338333
R734 VGND.n423 VGND.n1 0.0338333
R735 VGND.n419 VGND.n1 0.0338333
R736 VGND.n419 VGND.n418 0.0338333
R737 VGND.n416 VGND.n7 0.0338333
R738 VGND.n412 VGND.n7 0.0338333
R739 VGND.n412 VGND.n411 0.0338333
R740 VGND.n411 VGND.n410 0.0338333
R741 VGND.n418 VGND.n417 0.0329074
R742 VGND.n424 VGND.n0 0.0305926
R743 VGND.n315 VGND.n285 0.0236481
R744 VGND.n322 VGND.n321 0.0148519
R745 VGND.n312 VGND.n285 0.0106852
R746 VGND.n424 VGND.n423 0.00374074
R747 VGND.n417 VGND.n416 0.00142593
R748 OUT.n0 OUT.t0 662.732
R749 OUT.n1 OUT.t2 219.184
R750 OUT.n0 OUT.t1 131.75
R751 OUT OUT.n1 3.97095
R752 OUT.n1 OUT.n0 1.1255
R753 IN.n0 IN.t0 416.05
R754 IN.n0 IN.t1 322.983
R755 IN IN.n0 4.71567
R756 VDDOUT.n2 VDDOUT.t1 663.173
R757 VDDOUT.n1 VDDOUT.t3 663.153
R758 VDDOUT.n0 VDDOUT.t0 483.637
R759 VDDOUT.n0 VDDOUT.t2 428.365
R760 VDDOUT.n1 VDDOUT.n0 379.416
R761 VDDOUT VDDOUT.n2 0.3385
R762 VDDOUT.n2 VDDOUT.n1 0.006125
C0 a_1778_346# VDDOUT 0.313758f
C1 VDDIN a_897_442# 0.167083f
C2 IN VDDIN 0.224671f
C3 VDDIN a_373_442# 0.480793f
C4 OUT a_373_442# 0.204639f
C5 VDDIN VDDOUT 0.153557f
C6 OUT VDDOUT 0.505491f
C7 a_373_442# a_897_442# 0.43646f
C8 IN a_373_442# 0.209079f
C9 VDDOUT a_897_442# 0.037759f
C10 a_373_442# VDDOUT 0.0691f
C11 OUT a_1778_346# 0.340274f
C12 a_1778_346# a_897_442# 0.115354f
C13 a_1778_346# a_373_442# 0.158653f
C14 OUT VGND 0.778369f
C15 IN VGND 0.70206f
C16 VDDOUT VGND 3.37132f
C17 VDDIN VGND 3.68719f
C18 a_1778_346# VGND 0.315222f
C19 a_897_442# VGND 0.791735f
C20 a_373_442# VGND 1.39777f
.ends

